library verilog;
use verilog.vl_types.all;
entity Sersum_V8_vlg_check_tst is
    port(
        ssum            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Sersum_V8_vlg_check_tst;
