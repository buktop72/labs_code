-- Copyright (C) 1991-2010 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 9.1 Build 350 03/24/2010 Service Pack 2 SJ Web Edition
-- Created on Thu Nov 03 11:28:41 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY lab11_automat IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        a : IN STD_LOGIC := '0';
        b : IN STD_LOGIC := '0';
        q : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END lab11_automat;

ARCHITECTURE BEHAVIOR OF lab11_automat IS
    TYPE type_fstate IS (state3,state0,state1,state2,state4,state5,state14,state7,state8,state6,state13,state10,state15,state11,state12,state9);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,a,b)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state5;
            q <= "0000";
        ELSE
            q <= "0000";
            CASE fstate IS
                WHEN state3 =>
                    reg_fstate <= state11;

                    q <= "0011";
                WHEN state0 =>
                    IF ((a = '1')) THEN
                        reg_fstate <= state3;
                    ELSIF (NOT((a = '1'))) THEN
                        reg_fstate <= state14;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state0;
                    END IF;

                    q <= "0000";
                WHEN state1 =>
                    reg_fstate <= state9;

                    q <= "0001";
                WHEN state2 =>
                    reg_fstate <= state13;

                    q <= "0010";
                WHEN state4 =>
                    reg_fstate <= state2;

                    q <= "0100";
                WHEN state5 =>
                    reg_fstate <= state0;

                    q <= "0101";
                WHEN state14 =>
                    reg_fstate <= state8;

                    q <= "1110";
                WHEN state7 =>
                    IF (NOT((b = '1'))) THEN
                        reg_fstate <= state4;
                    ELSIF ((b = '1')) THEN
                        reg_fstate <= state6;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state7;
                    END IF;

                    q <= "0111";
                WHEN state8 =>
                    reg_fstate <= state7;

                    q <= "1000";
                WHEN state6 =>
                    reg_fstate <= state2;

                    q <= "0110";
                WHEN state13 =>
                    reg_fstate <= state10;

                    q <= "1101";
                WHEN state10 =>
                    reg_fstate <= state15;

                    q <= "1010";
                WHEN state15 =>
                    reg_fstate <= state5;

                    q <= "1111";
                WHEN state11 =>
                    IF ((b = '1')) THEN
                        reg_fstate <= state1;
                    ELSIF (NOT((b = '1'))) THEN
                        reg_fstate <= state12;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state11;
                    END IF;

                    q <= "1011";
                WHEN state12 =>
                    reg_fstate <= state9;

                    q <= "1100";
                WHEN state9 =>
                    reg_fstate <= state2;

                    q <= "1001";
                WHEN OTHERS => 
                    q <= "XXXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
