library verilog;
use verilog.vl_types.all;
entity Sersum_V8_vlg_vec_tst is
end Sersum_V8_vlg_vec_tst;
