library verilog;
use verilog.vl_types.all;
entity laba5 is
    port(
        y               : out    vl_logic;
        a1              : in     vl_logic;
        a0              : in     vl_logic;
        a2              : in     vl_logic
    );
end laba5;
