library verilog;
use verilog.vl_types.all;
entity laba5_vlg_check_tst is
    port(
        y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end laba5_vlg_check_tst;
