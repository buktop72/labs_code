// Copyright (C) 1991-2010 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 9.1 Build 350 03/24/2010 Service Pack 2 SJ Web Edition
// Created on Thu Nov 03 11:53:03 2022

// synthesis message_off 10175

`timescale 1ns/1ns

module lab11_automat (
    reset,clk,a,b,
    q[3:0]);

    input reset;
    input clk;
    input a;
    input b;
    tri0 reset;
    tri0 a;
    tri0 b;
    output [3:0] q;
    reg [3:0] q;
    reg [15:0] fstate;
    reg [15:0] reg_fstate;
    parameter state3=0,state0=1,state1=2,state2=3,state4=4,state5=5,state14=6,state7=7,state8=8,state6=9,state13=10,state10=11,state15=12,state11=13,state12=14,state9=15;

    always @(posedge clk)
    begin
        if (clk) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or a or b)
    begin
        if (reset) begin
            reg_fstate <= state5;
            q <= 4'b0000;
        end
        else begin
            q <= 4'b0000;
            case (fstate)
                state3: begin
                    reg_fstate <= state11;

                    q <= 4'b0011;
                end
                state0: begin
                    if (a)
                        reg_fstate <= state3;
                    else if (~(a))
                        reg_fstate <= state14;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state0;

                    q <= 4'b0000;
                end
                state1: begin
                    reg_fstate <= state9;

                    q <= 4'b0001;
                end
                state2: begin
                    reg_fstate <= state13;

                    q <= 4'b0010;
                end
                state4: begin
                    reg_fstate <= state2;

                    q <= 4'b0100;
                end
                state5: begin
                    reg_fstate <= state0;

                    q <= 4'b0101;
                end
                state14: begin
                    reg_fstate <= state8;

                    q <= 4'b1110;
                end
                state7: begin
                    if (~(b))
                        reg_fstate <= state4;
                    else if (b)
                        reg_fstate <= state6;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state7;

                    q <= 4'b0111;
                end
                state8: begin
                    reg_fstate <= state7;

                    q <= 4'b1000;
                end
                state6: begin
                    reg_fstate <= state2;

                    q <= 4'b0110;
                end
                state13: begin
                    reg_fstate <= state10;

                    q <= 4'b1101;
                end
                state10: begin
                    reg_fstate <= state15;

                    q <= 4'b1010;
                end
                state15: begin
                    reg_fstate <= state5;

                    q <= 4'b1111;
                end
                state11: begin
                    if (b)
                        reg_fstate <= state1;
                    else if (~(b))
                        reg_fstate <= state12;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state11;

                    q <= 4'b1011;
                end
                state12: begin
                    reg_fstate <= state9;

                    q <= 4'b1100;
                end
                state9: begin
                    reg_fstate <= state2;

                    q <= 4'b1001;
                end
                default: begin
                    q <= 4'bxxxx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // lab11_automat
