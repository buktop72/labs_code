library verilog;
use verilog.vl_types.all;
entity laba5_vlg_vec_tst is
end laba5_vlg_vec_tst;
